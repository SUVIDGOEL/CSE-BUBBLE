`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.04.2025 04:22:39
// Design Name: 
// Module Name: instruction_decode
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module instruction_decode(
    input [31:0] instruction,
    output [5:0] opcode,
    output [4:0] rs,
    output [4:0] rt,
    output [4:0] rd,
    output [4:0] shamt,
    output [6:0] funct,
    output [15:0] immediate,
    output [25:0] jump_target
);
    assign opcode = instruction [31:26];
    assign rs = instruction [25:21];
    assign rt = instruction [20:16];
    assign rd = instruction [15:11];
    assign shamt = instruction [10:6];
    assign funct = instruction [5:0];
    assign immediate = instruction [15:0];
    assign jump_target = instruction [25:0];  
endmodule